module demask(
    input clk,
    input srstn,
    input start,
    input [624:0] in,
    output reg finish,
    output reg [223:0] demask_out
);

parameter IDLE = 1'b0, OUT = 1'b1;

reg state, state_nxt;
reg [624:0] pattern, pattern_nxt;
reg [2:0] label;

always @(posedge clk) begin
    if(~srstn) state <= IDLE;
    else state <= state_nxt;
    pattern <= pattern_nxt;
end

always @(*) begin
    case(state) //synopsys parallel_case
    IDLE: state_nxt= (start) ? OUT : IDLE;
    OUT: state_nxt = IDLE;
    default: state_nxt = IDLE;
    endcase
end

always @(*) begin
    pattern_nxt = (start) ? in : pattern;
    label = {~pattern[422], pattern[421], ~pattern[420]};
    finish = (state) ? 1 : 0;
end

always @(*) begin
    case(label) //synopsys parallel_case
    3'b000: demask_out = {~pattern[0], pattern[1], pattern[25], ~pattern[26], ~pattern[50], pattern[51], pattern[75], ~pattern[76],
                          ~pattern[100], pattern[101], pattern[125], ~pattern[126], ~pattern[150], pattern[151], pattern[175], ~pattern[176],
                          ~pattern[200], pattern[201], pattern[225], ~pattern[226], ~pattern[250], pattern[251], pattern[275], ~pattern[276],
                          ~pattern[300], pattern[301], pattern[325], ~pattern[326], ~pattern[350], pattern[351], pattern[375], ~pattern[376],
                          pattern[377], ~pattern[378], ~pattern[352], pattern[353], pattern[327], ~pattern[328], ~pattern[302], pattern[303],
                          pattern[277], ~pattern[278], ~pattern[252], pattern[253], pattern[227], ~pattern[228], ~pattern[202], pattern[203],
                          pattern[177], ~pattern[178], ~pattern[152], pattern[153], pattern[127], ~pattern[128], ~pattern[102], pattern[103],
                          pattern[77],  ~pattern[78],  ~pattern[52],  pattern[53],  pattern[27],  ~pattern[28],  ~pattern[2],   pattern[3],
                          ~pattern[4], pattern[5], pattern[29], ~pattern[30], ~pattern[54], pattern[55], pattern[79], ~pattern[80],
                          pattern[229], ~pattern[230], ~pattern[254], pattern[255], pattern[279], ~pattern[280], ~pattern[304], pattern[305],
                          pattern[329], ~pattern[330], ~pattern[354], pattern[355], pattern[379], ~pattern[380], pattern[381], ~pattern[382],
                          ~pattern[356], pattern[357], pattern[331], ~pattern[332], ~pattern[306], pattern[307], pattern[281], ~pattern[282],
                          ~pattern[256], pattern[257], pattern[231], ~pattern[232], pattern[81], ~pattern[82], ~pattern[56], pattern[57],
                          pattern[31], ~pattern[32], ~pattern[6], pattern[7], ~pattern[8], pattern[9], pattern[33], ~pattern[34],
                          ~pattern[58], pattern[59], pattern[83], ~pattern[84], pattern[109], ~pattern[134], pattern[159], ~pattern[184],
                          pattern[209], pattern[233], ~pattern[234], ~pattern[258], pattern[259], pattern[283], ~pattern[284], ~pattern[308],
                          pattern[309], pattern[333], ~pattern[334], ~pattern[358], pattern[359], pattern[383], ~pattern[384], ~pattern[408],
                          pattern[409], pattern[433], ~pattern[434], pattern[483], ~pattern[484], ~pattern[508], pattern[509], pattern[533],
                          pattern[534], ~pattern[558], pattern[559], pattern[583], ~pattern[584], ~pattern[608], pattern[609], ~pattern[610],
                          pattern[611], pattern[585], ~pattern[586], ~pattern[560], pattern[561], pattern[535], ~pattern[536], ~pattern[510],
                          pattern[511], pattern[485], ~pattern[486], pattern[435], ~pattern[436], ~pattern[410], pattern[411], pattern[385],
                          ~pattern[386], ~pattern[360], pattern[361], pattern[335], ~pattern[336], ~pattern[310], pattern[311], pattern[285],
                          ~pattern[286], ~pattern[260], pattern[261], pattern[235], ~pattern[236], ~pattern[210], pattern[211], pattern[185],
                          ~pattern[186], ~pattern[160], pattern[161], pattern[135], ~pattern[136], ~pattern[110], pattern[111], pattern[85],
                          ~pattern[86], ~pattern[60], pattern[61], pattern[35], ~pattern[36], ~pattern[10], pattern[11], ~pattern[12],
                          pattern[13], pattern[37], ~pattern[38], ~pattern[62], pattern[63], pattern[87], ~pattern[88], ~pattern[112],
                          pattern[113], pattern[137], ~pattern[138], ~pattern[162], pattern[163], pattern[187], ~pattern[188], ~pattern[212],
                          pattern[213], pattern[237], ~pattern[238], ~pattern[262], pattern[263], pattern[287], ~pattern[288], ~pattern[312]};

    3'b001: demask_out = {~pattern[0], ~pattern[1], pattern[25], pattern[26], ~pattern[50], ~pattern[51], pattern[75], pattern[76],
                          ~pattern[100], ~pattern[101], pattern[125], pattern[126], ~pattern[150], ~pattern[151], pattern[175], pattern[176],
                          ~pattern[200], ~pattern[201], pattern[225], pattern[226], ~pattern[250], ~pattern[251], pattern[275], pattern[276],
                          ~pattern[300], ~pattern[301], pattern[325], pattern[326], ~pattern[350], ~pattern[351], pattern[375], pattern[376],
                          pattern[377], pattern[378], ~pattern[352], ~pattern[353], pattern[327], pattern[328], ~pattern[302], ~pattern[303],
                          pattern[277], pattern[278], ~pattern[252], ~pattern[253], pattern[227], pattern[228], ~pattern[202], ~pattern[203],
                          pattern[177], pattern[178], ~pattern[152], ~pattern[153], pattern[127], pattern[128], ~pattern[102], ~pattern[103],
                          pattern[77],  pattern[78],  ~pattern[52],  ~pattern[53],  pattern[27],  pattern[28],  ~pattern[2],   ~pattern[3],
                          ~pattern[4], ~pattern[5], pattern[29], pattern[30], ~pattern[54], ~pattern[55], pattern[79], pattern[80],
                          pattern[229], pattern[230], ~pattern[254], ~pattern[255], pattern[279], pattern[280], ~pattern[304], ~pattern[305],
                          pattern[329], pattern[330], ~pattern[354], ~pattern[355], pattern[379], pattern[380], pattern[381], pattern[382],
                          ~pattern[356], ~pattern[357], pattern[331], pattern[332], ~pattern[306], ~pattern[307], pattern[281], pattern[282],
                          ~pattern[256], ~pattern[257], pattern[231], pattern[232], pattern[81], pattern[82], ~pattern[56], ~pattern[57],
                          pattern[31], pattern[32], ~pattern[6], ~pattern[7], ~pattern[8], ~pattern[9], pattern[33], pattern[34],
                          ~pattern[58], ~pattern[59], pattern[83], pattern[84], ~pattern[109], pattern[134], ~pattern[159], pattern[184],
                          ~pattern[209], pattern[233], pattern[234], ~pattern[258], ~pattern[259], pattern[283], pattern[284], ~pattern[308],
                          ~pattern[309], pattern[333], pattern[334], ~pattern[358], ~pattern[359], pattern[383], pattern[384], ~pattern[408],
                          ~pattern[409], pattern[433], pattern[434], pattern[483], pattern[484], ~pattern[508], ~pattern[509], pattern[533],
                          pattern[534], ~pattern[558], ~pattern[559], pattern[583], pattern[584], ~pattern[608], ~pattern[609], ~pattern[610],
                          ~pattern[611], pattern[585], pattern[586], ~pattern[560], ~pattern[561], pattern[535], pattern[536], ~pattern[510],
                          ~pattern[511], pattern[485], pattern[486], pattern[435], pattern[436], ~pattern[410], ~pattern[411], pattern[385],
                          pattern[386], ~pattern[360], ~pattern[361], pattern[335], pattern[336], ~pattern[310], ~pattern[311], pattern[285],
                          pattern[286], ~pattern[260], ~pattern[261], pattern[235], pattern[236], ~pattern[210], ~pattern[211], pattern[185],
                          pattern[186], ~pattern[160], ~pattern[161], pattern[135], pattern[136], ~pattern[110], ~pattern[111], pattern[85],
                          pattern[86], ~pattern[60], ~pattern[61], pattern[35], pattern[36], ~pattern[10], ~pattern[11], ~pattern[12],
                          ~pattern[13], pattern[37], pattern[38], ~pattern[62], ~pattern[63], pattern[87], pattern[88], ~pattern[112],
                          ~pattern[113], pattern[137], pattern[138], ~pattern[162], ~pattern[163], pattern[187], pattern[188], ~pattern[212],
                          ~pattern[213], pattern[237], pattern[238], ~pattern[262], ~pattern[263], pattern[287], pattern[288], ~pattern[312]};

    3'b010: demask_out = {~pattern[0],   pattern[1],   ~pattern[25],  pattern[26],  ~pattern[50],  pattern[51],  ~pattern[75],  pattern[76],
                          ~pattern[100], pattern[101], ~pattern[125], pattern[126], ~pattern[150], pattern[151], ~pattern[175], pattern[176],
                          ~pattern[200], pattern[201], ~pattern[225], pattern[226], ~pattern[250], pattern[251], ~pattern[275], pattern[276],
                          ~pattern[300], pattern[301], ~pattern[325], pattern[326], ~pattern[350], pattern[351], ~pattern[375], pattern[376],
                          pattern[377], ~pattern[378], pattern[352], ~pattern[353], pattern[327], ~pattern[328], pattern[302], ~pattern[303],
                          pattern[277], ~pattern[278], pattern[252], ~pattern[253], pattern[227], ~pattern[228], pattern[202], ~pattern[203],
                          pattern[177], ~pattern[178], pattern[152], ~pattern[153], pattern[127], ~pattern[128], pattern[102], ~pattern[103],
                          pattern[77],  ~pattern[78],  pattern[52],  ~pattern[53],  pattern[27],  ~pattern[28],  pattern[2],   ~pattern[3],
                          pattern[4],   pattern[5],   pattern[29],  pattern[30],  pattern[54],  pattern[55],  pattern[79],  pattern[80],
                          pattern[229], pattern[230], pattern[254], pattern[255], pattern[279], pattern[280], pattern[304], pattern[305],
                          pattern[329], pattern[330], pattern[354], pattern[355], pattern[379], pattern[380], ~pattern[381], pattern[382],
                          ~pattern[356], pattern[357], ~pattern[331], pattern[332], ~pattern[306], pattern[307], ~pattern[281], pattern[282],
                          ~pattern[256], pattern[257], ~pattern[231], pattern[232], ~pattern[81],  pattern[82],  ~pattern[56],  pattern[57],
                          ~pattern[31],  pattern[32],  ~pattern[6],   pattern[7],   pattern[8],   ~pattern[9],   pattern[33],  ~pattern[34],
                          pattern[58],  ~pattern[59],  pattern[83],  ~pattern[84],  ~pattern[109], ~pattern[134], ~pattern[159], ~pattern[184],
                          ~pattern[209], pattern[233], ~pattern[234], pattern[258], ~pattern[259], pattern[283], ~pattern[284], pattern[308],
                          ~pattern[309], pattern[333], ~pattern[334], pattern[358], ~pattern[359], pattern[383], ~pattern[384], pattern[408],
                          ~pattern[409], pattern[433],~pattern[434], pattern[483], ~pattern[484], pattern[508], ~pattern[509], pattern[533],
                          ~pattern[534], pattern[558], ~pattern[559], pattern[583], ~pattern[584], pattern[608], ~pattern[609], pattern[610],
                          pattern[611], pattern[585], pattern[586], pattern[560], pattern[561], pattern[535], pattern[536], pattern[510],
                          pattern[511], pattern[485], pattern[486], pattern[435], pattern[436], pattern[410], pattern[411], pattern[385],
                          pattern[386], pattern[360], pattern[361], pattern[335], pattern[336], pattern[310], pattern[311], pattern[285],
                          pattern[286], pattern[260], pattern[261], pattern[235], pattern[236], pattern[210], pattern[211], pattern[185],
                          pattern[186], pattern[160], pattern[161], pattern[135], pattern[136], pattern[110], pattern[111], pattern[85],
                          pattern[86],  pattern[60],  pattern[61],  pattern[35],  pattern[36],  pattern[10],  pattern[11],  ~pattern[12],
                          pattern[13],  ~pattern[37],  pattern[38],  ~pattern[62],  pattern[63],  ~pattern[87],  pattern[88],  ~pattern[112],
                          pattern[113], ~pattern[137], pattern[138], ~pattern[162], pattern[163], ~pattern[187], pattern[188], ~pattern[212],
                          pattern[213], ~pattern[237], pattern[238], ~pattern[262], pattern[263],~pattern[287], pattern[288], ~pattern[312]};

    3'b011: demask_out = {~pattern[0],   pattern[1],   pattern[25],  pattern[26],  pattern[50], ~pattern[51], ~pattern[75],  pattern[76],
                          pattern[100], pattern[101], pattern[125], ~pattern[126], ~pattern[150], pattern[151], pattern[175], pattern[176],
                          pattern[200], ~pattern[201], ~pattern[225], pattern[226], pattern[250], pattern[251], pattern[275], ~pattern[276],
                          ~pattern[300], pattern[301], pattern[325], pattern[326], pattern[350], ~pattern[351], ~pattern[375], pattern[376],
                          pattern[377], ~pattern[378], pattern[352], pattern[353], ~pattern[327], pattern[328], pattern[302], ~pattern[303],
                          pattern[277], pattern[278], ~pattern[252], pattern[253], pattern[227], ~pattern[228], pattern[202], pattern[203],
                          ~pattern[177], pattern[178], pattern[152], ~pattern[153], pattern[127], pattern[128], ~pattern[102], pattern[103],
                          pattern[77],  ~pattern[78],  pattern[52],  pattern[53],  ~pattern[27],  pattern[28],  pattern[2],   ~pattern[3],
                          pattern[4],   pattern[5],   pattern[29],  ~pattern[30], ~pattern[54],  pattern[55],  pattern[79],  pattern[80],
                          pattern[229], pattern[230], pattern[254], ~pattern[255], ~pattern[279], pattern[280], pattern[304], pattern[305],
                          pattern[329], ~pattern[330], ~pattern[354], pattern[355], pattern[379], pattern[380], ~pattern[381], pattern[382],
                          pattern[356], ~pattern[357], pattern[331], pattern[332], ~pattern[306], pattern[307], pattern[281], ~pattern[282],
                          pattern[256], pattern[257], ~pattern[231], pattern[232], ~pattern[81],  pattern[82],  pattern[56],  ~pattern[57],
                          pattern[31],  pattern[32],  ~pattern[6],   pattern[7],   pattern[8],  ~pattern[9],  ~pattern[33],  pattern[34],
                          pattern[58],  pattern[59],  pattern[83],  ~pattern[84],  pattern[109], pattern[134], ~pattern[159], pattern[184],
                          pattern[209], pattern[233], ~pattern[234], ~pattern[258], pattern[259], pattern[283], pattern[284], pattern[308],
                          ~pattern[309], ~pattern[333], pattern[334], pattern[358], pattern[359], pattern[383], ~pattern[384], ~pattern[408],
                          pattern[409], pattern[433], pattern[434], ~pattern[483], pattern[484], pattern[508], pattern[509], pattern[533],
                          pattern[534], pattern[558], pattern[559], pattern[583], pattern[584], pattern[608], ~pattern[609], pattern[610],
                          pattern[611], ~pattern[585], pattern[586], pattern[560], pattern[561], pattern[535], pattern[536], ~pattern[510],
                          pattern[511], pattern[485], ~pattern[486], ~pattern[435], pattern[436], pattern[410], ~pattern[411], pattern[385],
                          pattern[386], ~pattern[360], pattern[361], pattern[335], ~pattern[336], pattern[310], pattern[311], ~pattern[285],
                          pattern[286], pattern[260], ~pattern[261], pattern[235], pattern[236], ~pattern[210], pattern[211], pattern[185],
                          ~pattern[186], pattern[160], pattern[161], ~pattern[135], pattern[136], pattern[110], ~pattern[111], pattern[85],
                          pattern[86],  ~pattern[60],  pattern[61],  pattern[35],  ~pattern[36],  pattern[10],  pattern[11],  ~pattern[12],
                          pattern[13],  pattern[37],  pattern[38],  pattern[62],  ~pattern[63], ~pattern[87],  pattern[88],  pattern[112],
                          pattern[113], pattern[137], ~pattern[138], ~pattern[162], pattern[163], pattern[187], pattern[188], pattern[212],
                          ~pattern[213], ~pattern[237], pattern[238], pattern[262], pattern[263], pattern[287], ~pattern[288], ~pattern[312]};

    3'b100: demask_out = {~pattern[0],   pattern[1],   pattern[25],  ~pattern[26],  pattern[50],  ~pattern[51],  ~pattern[75],  pattern[76],
                          ~pattern[100], pattern[101], pattern[125], ~pattern[126], pattern[150], ~pattern[151], ~pattern[175], pattern[176],
                          ~pattern[200], pattern[201], pattern[225], ~pattern[226], pattern[250], ~pattern[251], ~pattern[275], pattern[276],
                          ~pattern[300], pattern[301], pattern[325], ~pattern[326], pattern[350], ~pattern[351], ~pattern[375], pattern[376],
                          pattern[377], pattern[378], ~pattern[352], ~pattern[353], ~pattern[327], ~pattern[328], pattern[302], pattern[303],
                          pattern[277], pattern[278], ~pattern[252], ~pattern[253], ~pattern[227], ~pattern[228], pattern[202], pattern[203],
                          pattern[177], pattern[178], ~pattern[152], ~pattern[153], ~pattern[127], ~pattern[128], pattern[102], pattern[103],
                          pattern[77],  pattern[78],  ~pattern[52],  ~pattern[53],  ~pattern[27],  ~pattern[28],  pattern[2],   pattern[3],
                          ~pattern[4],   ~pattern[5],   pattern[29],  pattern[30],  pattern[54],  pattern[55],  ~pattern[79],  ~pattern[80],
                          pattern[229], pattern[230], pattern[254], pattern[255], ~pattern[279], ~pattern[280], ~pattern[304], ~pattern[305],
                          pattern[329], pattern[330], pattern[354], pattern[355], ~pattern[379], ~pattern[380], ~pattern[381], pattern[382],
                          pattern[356], ~pattern[357], pattern[331], ~pattern[332], ~pattern[306], pattern[307], ~pattern[281], pattern[282],
                          pattern[256], ~pattern[257], pattern[231], ~pattern[232], ~pattern[81],  pattern[82],  pattern[56],  ~pattern[57],
                          pattern[31],  ~pattern[32],  ~pattern[6],   pattern[7],   pattern[8],   pattern[9],   ~pattern[33],  ~pattern[34],
                          ~pattern[58],  ~pattern[59],  pattern[83],  pattern[84],  pattern[109], ~pattern[134], ~pattern[159], pattern[184],
                          pattern[209], ~pattern[233], ~pattern[234], ~pattern[258], ~pattern[259], pattern[283], pattern[284], pattern[308],
                          pattern[309], ~pattern[333], ~pattern[334], ~pattern[358], ~pattern[359], pattern[383], pattern[384], pattern[408],
                          pattern[409], ~pattern[433], ~pattern[434], pattern[483], pattern[484], pattern[508], pattern[509], ~pattern[533],
                          ~pattern[534], ~pattern[558], ~pattern[559], pattern[583], pattern[584], pattern[608], pattern[609], ~pattern[610],
                          ~pattern[611], ~pattern[585], ~pattern[586], pattern[560], pattern[561], pattern[535], pattern[536], ~pattern[510],
                          ~pattern[511], ~pattern[485], ~pattern[486], pattern[435], pattern[436], ~pattern[410], ~pattern[411], ~pattern[385],
                          ~pattern[386], pattern[360], pattern[361], pattern[335], pattern[336], ~pattern[310], ~pattern[311], ~pattern[285],
                          ~pattern[286], pattern[260], pattern[261], pattern[235], pattern[236], ~pattern[210], ~pattern[211], ~pattern[185],
                          ~pattern[186], pattern[160], pattern[161], pattern[135], pattern[136], ~pattern[110], ~pattern[111], ~pattern[85],
                          ~pattern[86],  pattern[60],  pattern[61],  pattern[35],  pattern[36],  ~pattern[10],  ~pattern[11],  ~pattern[12],
                          pattern[13],  pattern[37],  ~pattern[38],  pattern[62],  ~pattern[63],  ~pattern[87],  pattern[88],  ~pattern[112],
                          pattern[113], pattern[137], ~pattern[138], pattern[162], ~pattern[163], ~pattern[187], pattern[188], ~pattern[212],
                          pattern[213], pattern[237], ~pattern[238], pattern[262], ~pattern[263], ~pattern[287], pattern[288], ~pattern[312]};

    3'b101: demask_out = {~pattern[0],   ~pattern[1],   ~pattern[25],  pattern[26],  ~pattern[50],  pattern[51],  ~pattern[75],  pattern[76],
                          ~pattern[100], pattern[101], ~pattern[125], pattern[126], ~pattern[150], ~pattern[151], ~pattern[175], pattern[176],
                          ~pattern[200], pattern[201], ~pattern[225], pattern[226], ~pattern[250], pattern[251], ~pattern[275], pattern[276],
                          ~pattern[300], ~pattern[301], ~pattern[325], pattern[326], ~pattern[350], pattern[351], ~pattern[375], pattern[376],
                          ~pattern[377], pattern[378], pattern[352], ~pattern[353], pattern[327], pattern[328], ~pattern[302], ~pattern[303],
                          pattern[277], pattern[278], pattern[252], ~pattern[253], ~pattern[227], pattern[228], pattern[202], ~pattern[203],
                          pattern[177], pattern[178], ~pattern[152], ~pattern[153], pattern[127], pattern[128], pattern[102], ~pattern[103],
                          ~pattern[77],  pattern[78],  pattern[52],  ~pattern[53],  pattern[27],  pattern[28],  ~pattern[2],   ~pattern[3],
                          ~pattern[4],   ~pattern[5],   pattern[29],  pattern[30],  pattern[54],  pattern[55],  ~pattern[79],  pattern[80],
                          ~pattern[229], pattern[230], pattern[254], pattern[255], pattern[279], pattern[280], ~pattern[304], ~pattern[305],
                          pattern[329], pattern[330], pattern[354], pattern[355], ~pattern[379], pattern[380], ~pattern[381], pattern[382],
                          ~pattern[356], pattern[357], ~pattern[331], pattern[332], ~pattern[306], ~pattern[307], ~pattern[281], pattern[282],
                          ~pattern[256], pattern[257], ~pattern[231], pattern[232], ~pattern[81],  pattern[82],  ~pattern[56],  pattern[57],
                          ~pattern[31],  pattern[32],  ~pattern[6],   ~pattern[7],   ~pattern[8],   ~pattern[9],   pattern[33],  pattern[34],
                          pattern[58],  ~pattern[59],  ~pattern[83],  pattern[84],  ~pattern[109], pattern[134], ~pattern[159], pattern[184],
                          ~pattern[209], ~pattern[233], pattern[234], pattern[258], ~pattern[259], pattern[283], pattern[284], ~pattern[308],
                          ~pattern[309], pattern[333], pattern[334], pattern[358], ~pattern[359], ~pattern[383], pattern[384], pattern[408],
                          ~pattern[409], pattern[433], pattern[434], pattern[483], pattern[484], pattern[508], ~pattern[509], ~pattern[533],
                          pattern[534], pattern[558], ~pattern[559], pattern[583], pattern[584], ~pattern[608], ~pattern[609], ~pattern[610],
                          ~pattern[611], pattern[585], pattern[586], pattern[560], pattern[561], ~pattern[535], pattern[536], pattern[510],
                          pattern[511], pattern[485], pattern[486], pattern[435], pattern[436], pattern[410], pattern[411], ~pattern[385],
                          pattern[386], pattern[360], pattern[361], pattern[335], pattern[336], ~pattern[310], ~pattern[311], pattern[285],
                          pattern[286], pattern[260], pattern[261], ~pattern[235], pattern[236], pattern[210], pattern[211], pattern[185],
                          pattern[186], ~pattern[160], ~pattern[161], pattern[135], pattern[136], pattern[110], pattern[111], ~pattern[85],
                          pattern[86],  pattern[60],  pattern[61],  pattern[35],  pattern[36],  ~pattern[10],  ~pattern[11],  ~pattern[12],
                          ~pattern[13],  ~pattern[37],  pattern[38],  ~pattern[62],  pattern[63],  ~pattern[87],  pattern[88],  ~pattern[112],
                          pattern[113], ~pattern[137], pattern[138], ~pattern[162], ~pattern[163], ~pattern[187], pattern[188], ~pattern[212],
                          pattern[213], ~pattern[237], pattern[238], ~pattern[262], pattern[263], ~pattern[287], pattern[288], ~pattern[312]};

    3'b110: demask_out = {~pattern[0],   ~pattern[1],   ~pattern[25],  ~pattern[26],  ~pattern[50],  ~pattern[51],  ~pattern[75],  pattern[76],
                          ~pattern[100], pattern[101], ~pattern[125], pattern[126], ~pattern[150], ~pattern[151], ~pattern[175], ~pattern[176],
                          ~pattern[200], ~pattern[201], ~pattern[225], pattern[226], ~pattern[250], pattern[251], ~pattern[275], pattern[276],
                          ~pattern[300], ~pattern[301], ~pattern[325], ~pattern[326], ~pattern[350], ~pattern[351], ~pattern[375], pattern[376],
                          ~pattern[377], pattern[378], pattern[352], ~pattern[353], ~pattern[327], pattern[328], ~pattern[302], ~pattern[303],
                          pattern[277], pattern[278], ~pattern[252], ~pattern[253], ~pattern[227], pattern[228], pattern[202], ~pattern[203],
                          ~pattern[177], pattern[178], ~pattern[152], ~pattern[153], pattern[127], pattern[128], ~pattern[102], ~pattern[103],
                          ~pattern[77],  pattern[78],  pattern[52],  ~pattern[53],  ~pattern[27],  pattern[28],  ~pattern[2],   ~pattern[3],
                          ~pattern[4],   ~pattern[5],   pattern[29],  pattern[30],  ~pattern[54],  pattern[55],  ~pattern[79],  pattern[80],
                          ~pattern[229], pattern[230], pattern[254], ~pattern[255], ~pattern[279], ~pattern[280], ~pattern[304], ~pattern[305],
                          pattern[329], pattern[330], ~pattern[354], pattern[355], ~pattern[379], pattern[380], ~pattern[381], pattern[382],
                          ~pattern[356], ~pattern[357], ~pattern[331], ~pattern[332], ~pattern[306], ~pattern[307], ~pattern[281], pattern[282],
                          ~pattern[256], pattern[257], ~pattern[231], pattern[232], ~pattern[81],  pattern[82],  ~pattern[56],  ~pattern[57],
                          ~pattern[31],  ~pattern[32],  ~pattern[6],   ~pattern[7],   ~pattern[8],   ~pattern[9],   ~pattern[33],  pattern[34],
                          pattern[58],  ~pattern[59],  ~pattern[83],  pattern[84],  ~pattern[109], pattern[134], ~pattern[159], pattern[184],
                          ~pattern[209], ~pattern[233], pattern[234], ~pattern[258], ~pattern[259], pattern[283], pattern[284], ~pattern[308],
                          ~pattern[309], ~pattern[333], pattern[334], pattern[358], ~pattern[359], ~pattern[383], pattern[384], ~pattern[408],
                          ~pattern[409], pattern[433], pattern[434], ~pattern[483], pattern[484], pattern[508], ~pattern[509], ~pattern[533],
                          pattern[534], ~pattern[558], ~pattern[559], pattern[583], pattern[584], ~pattern[608], ~pattern[609], ~pattern[610],
                          ~pattern[611], ~pattern[585], ~pattern[586], pattern[560], ~pattern[561], ~pattern[535], pattern[536], ~pattern[510],
                          pattern[511], pattern[485], pattern[486], ~pattern[435], ~pattern[436], pattern[410], ~pattern[411], ~pattern[385],
                          pattern[386], ~pattern[360], pattern[361], pattern[335], pattern[336], ~pattern[310], ~pattern[311], ~pattern[285],
                          ~pattern[286], pattern[260], ~pattern[261], ~pattern[235], pattern[236], ~pattern[210], pattern[211], pattern[185],
                          pattern[186], ~pattern[160], ~pattern[161], ~pattern[135], ~pattern[136], pattern[110], ~pattern[111], ~pattern[85],
                          pattern[86],  ~pattern[60],  pattern[61],  pattern[35],  pattern[36],  ~pattern[10],  ~pattern[11],  ~pattern[12],
                          ~pattern[13],  ~pattern[37],  ~pattern[38],  ~pattern[62],  ~pattern[63],  ~pattern[87],  pattern[88],  ~pattern[112],
                          pattern[113], ~pattern[137], pattern[138], ~pattern[162], ~pattern[163], ~pattern[187], ~pattern[188], ~pattern[212],
                          ~pattern[213], ~pattern[237], pattern[238], ~pattern[262], pattern[263], ~pattern[287], pattern[288], ~pattern[312]};

    3'b111: demask_out = {~pattern[0],   pattern[1],   pattern[25],  pattern[26],  ~pattern[50],  pattern[51],  pattern[75],  ~pattern[76],
                          ~pattern[100], ~pattern[101], pattern[125], ~pattern[126], ~pattern[150], pattern[151], pattern[175], pattern[176],
                          ~pattern[200], pattern[201], pattern[225], ~pattern[226], ~pattern[250], ~pattern[251], pattern[275], ~pattern[276],
                          ~pattern[300], pattern[301], pattern[325], pattern[326], ~pattern[350], pattern[351], pattern[375], ~pattern[376],
                          pattern[377], ~pattern[378], pattern[352], pattern[353], pattern[327], ~pattern[328], ~pattern[302], pattern[303],
                          ~pattern[277], ~pattern[278], ~pattern[252], pattern[253], pattern[227], ~pattern[228], pattern[202], pattern[203],
                          pattern[177], ~pattern[178], ~pattern[152], pattern[153], ~pattern[127], ~pattern[128], ~pattern[102], pattern[103],
                          pattern[77],  ~pattern[78],  pattern[52],  pattern[53],  pattern[27],  ~pattern[28],  ~pattern[2],   pattern[3],
                          ~pattern[4],   pattern[5],   ~pattern[29],  ~pattern[30],  ~pattern[54],  ~pattern[55],  pattern[79],  ~pattern[80],
                          pattern[229], ~pattern[230], pattern[254], pattern[255], pattern[279], pattern[280], ~pattern[304], pattern[305],
                          ~pattern[329], ~pattern[330], ~pattern[354], ~pattern[355], pattern[379], ~pattern[380], pattern[381], ~pattern[382],
                          ~pattern[356], pattern[357], pattern[331], pattern[332], ~pattern[306], pattern[307], pattern[281], ~pattern[282],
                          ~pattern[256], ~pattern[257], pattern[231], ~pattern[232], pattern[81],  ~pattern[82],  ~pattern[56],  pattern[57],
                          pattern[31],  pattern[32],  ~pattern[6],   pattern[7],   ~pattern[8],   pattern[9],   pattern[33],  ~pattern[34],
                          pattern[58],  pattern[59],  pattern[83],  ~pattern[84],  pattern[109], ~pattern[134], pattern[159], ~pattern[184],
                          pattern[209], pattern[233], ~pattern[234], ~pattern[258], pattern[259], ~pattern[283], ~pattern[284], ~pattern[308],
                          pattern[309], pattern[333], ~pattern[334], pattern[358], pattern[359], pattern[383], ~pattern[384], ~pattern[408],
                          pattern[409], ~pattern[433], ~pattern[434], pattern[483], ~pattern[484], pattern[508], pattern[509], pattern[533],
                          ~pattern[534], ~pattern[558], pattern[559], ~pattern[583], ~pattern[584], ~pattern[608], pattern[609], ~pattern[610],
                          pattern[611], pattern[585], pattern[586], pattern[560], pattern[561], pattern[535], ~pattern[536], ~pattern[510],
                          ~pattern[511], ~pattern[485], ~pattern[486], pattern[435], pattern[436], pattern[410], pattern[411], pattern[385],
                          ~pattern[386], ~pattern[360], ~pattern[361], ~pattern[335], ~pattern[336], ~pattern[310], pattern[311], pattern[285],
                          pattern[286], pattern[260], pattern[261], pattern[235], ~pattern[236], ~pattern[210], ~pattern[211], ~pattern[185],
                          ~pattern[186], ~pattern[160], pattern[161], pattern[135], pattern[136], pattern[110], pattern[111], pattern[85],
                          ~pattern[86],  ~pattern[60],  ~pattern[61],  ~pattern[35],  ~pattern[36],  ~pattern[10],  pattern[11],  ~pattern[12],
                          pattern[13],  pattern[37],  pattern[38],  ~pattern[62],  pattern[63],  pattern[87],  ~pattern[88],  ~pattern[112],
                          ~pattern[113], pattern[137], ~pattern[138], ~pattern[162], pattern[163], pattern[187], pattern[188], ~pattern[212],
                          pattern[213], pattern[237], ~pattern[238], ~pattern[262], ~pattern[263], pattern[287], ~pattern[288], ~pattern[312]};     
    endcase
end

endmodule